library verilog;
use verilog.vl_types.all;
entity sobel_edge_tb is
end sobel_edge_tb;
